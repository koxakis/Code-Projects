module encoder(sel, res);

	input [7:0] res;
	
	output [2:0] sel;
	
	reg [7:0] sel;
	
	always @(res)
	begin
		case( sel)


endmodule 